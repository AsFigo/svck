# ----------------------------------------------------
# SPDX-FileCopyrightText: AsFigo Technologies, UK
# SPDX-FileCopyrightText: VerifWorks, India
# SPDX-License-Identifier: MIT
# ----------------------------------------------------

package p1;
  int tt;
endpackage

  int i1;

class c;
  rand int t;
  local int lvar_i1;
endclass : c

